module box(input [5:0] box_X,box_Y,
				 output logic [4:0] box_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h2, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1,
5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1, 5'h2, 5'h2, 5'h1, 5'h2, 5'h1, 5'h2, 5'h2, 5'h1, 5'h1,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h1,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2, 5'h2,
5'h3, 5'h2, 5'h2, 5'h2, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h2, 5'h2	};

	assign box_color_out = ROM[box_Y*40+box_X];


endmodule


module grass(input [5:0] grass_X,grass_Y,
				 output logic [4:0] grass_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5,
5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h4, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h6, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h5, 5'h4, 5'h4, 5'h4, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h4, 5'h4, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h6, 5'h6, 5'h6, 5'h6, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 5'h5, 
5'h5, 5'h5, 5'h4, 5'h4, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5, 5'h5, 5'h5, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h4, 5'h5};
	assign grass_color_out = ROM[grass_Y*40+grass_X];


endmodule


module brick(input [5:0] brick_X,brick_Y,
				 output logic [4:0] brick_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h8, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 5'h8, 5'h7, 5'h7, 5'h7, 5'h8, 5'h7, 5'h7, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h7, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 
5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h7, 5'h7, 5'h7, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h8, 5'h8, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 
5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9, 5'h9};
	assign brick_color_out = ROM[brick_Y*40+brick_X];


endmodule


module player(input [5:0] player_X,player_Y,
				 output logic [4:0] player_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hE, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'hE, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hD, 5'hD, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hD, 5'hD, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hD, 5'hD, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hD, 5'hD, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hD, 5'hD, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hD, 5'hD, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hD, 5'hD, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hD, 5'hD, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'hE, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'h1, 5'h1, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h1, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'h1, 5'h1, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'h1, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF};
	assign player_color_out = ROM[player_Y*40+player_X];


endmodule


module bomb( input [5:0] bomb_X,bomb_Y,
				 output logic [4:0] bomb_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hF, 5'hB, 5'hB, 5'hA, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 
5'hF, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 
5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hF, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hF, 5'hC, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hC, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 
5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 
5'hF, 5'hF, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 
5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hC, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hA, 5'hA, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hA, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hC, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF};
	assign bomb_color_out = ROM[bomb_Y*40+bomb_X];


endmodule

module explosion( input [5:0] explosion_X,explosion_Y,
				 output logic [4:0] explosion_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA};
	assign explosion_color_out = ROM[explosion_Y*40+explosion_X];


endmodule

//module heart();

module shoe( input [5:0] shoe_X,shoe_Y,
				 output logic [4:0] shoe_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hC, 5'hC, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h0, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'hC, 5'hC, 5'hC, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'h0, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'h0, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hC, 5'hB, 5'hC, 5'h0, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h8, 5'hB, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hC, 5'hC, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF};

	assign shoe_color_out = ROM[shoe_Y*40+shoe_X];
endmodule

module potion( input [5:0] potion_X,potion_Y,
				 output logic [4:0] potion_color_out
);
	parameter width = 40;
	parameter height = 40;
	parameter DATA_WIDTH = 5;
	parameter[0:height*width-1][DATA_WIDTH-1:0] ROM = {
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hC, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hC, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hB, 5'hB, 5'hC, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hC, 5'hA, 5'hA, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hE, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hE, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hC, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF};
	assign potion_color_out = ROM[potion_Y*40+potion_X];
endmodule